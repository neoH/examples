module top; // {
	cb_if t_if();
endmodule // }
